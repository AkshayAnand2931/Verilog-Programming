module tb;
    reg clk,clear,load,count;
    reg [2:0]i;
    wire cout;
    wire [2:0]o;
endmodule