module tb;
    reg a;
    reg b;
    wire c,d;
    and1 a1(a,b,c,d);

    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0,tb);
    end
    initial begin
        $monitor($time,a,b,c,d);
        a = 1'b0;
        b = 1'b0;
        #10
        a = 1'b0;
        b = 1'b1;
        #10
        a = 1'b1;
        b = 1'b0;
        #10
        a = 1'b1;
        b = 1'b1;
    end
endmodule